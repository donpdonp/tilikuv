module matrix

pub struct Message {
pub:
	room    string
	user    string
	message string
}
