module irc

pub struct Message {
pub:
	network string
	nick    string
	channel string
	message string
}
