module msg

struct IrcMsg {
}
