module msg

pub struct MatrixMsg {
}
