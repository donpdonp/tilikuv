module msg

pub struct IrcMsg {
}
