module msg

struct MatrixMsg {
}
